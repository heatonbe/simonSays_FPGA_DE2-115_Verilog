library verilog;
use verilog.vl_types.all;
entity simonSaysVGA_vlg_vec_tst is
end simonSaysVGA_vlg_vec_tst;
